----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:40:35 10/14/2023 
-- Design Name: 
-- Module Name:    desl_esq - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity desl_esq is                                           --Desloca todos os bits da entrada para a esquerda. Adiciona-se um '0' na posição mais à direita
    Port ( a : in  STD_LOGIC_VECTOR (3 downto 0);            --Entrada, o número binário de 4 bits do qual se quer fazer o deslocamento
           s : out  STD_LOGIC_VECTOR (3 downto 0);           --Resultado da operação, que retorna o delocamento à esquerda da entrada dada
	   bit_sinal : out STD_LOGIC;                        --Flag de sinal, apontando se o resultado da operação é positivo (0) ou negativo (1)
	   zero : out STD_LOGIC);                            --Flag de zero, apontando se o resultado da operação é o valor zero ("0000")
end desl_esq;

architecture Behavioral of desl_esq is

signal z : STD_LOGIC_VECTOR (3 downto 0);

begin

--Deslocamento dos bits: o bit da posição n recebe o bit da posição n-1. Como o bit mais à direita (bit 0) não possui um correspondente, receberá sempre 0
z(3) <= a(2);
z(2) <= a(1);
z(1) <= a(0);
z(0) <= '0';

s <= z;

bit_sinal <= a(2);               --O bit de sinal do resultado da operação de deslocamento à esquerda é z(3), que é equivalente a a(2) 

zero <= '1' when z = "0000" else '0';

end Behavioral;

